library ieee;
use ieee.STD_logic_1164.all;

entity MapeoLaberinto is
PORT ( 
		
		
		);


end MapeoLaberinto;

architecture behave of MapeoLaberinto is

begin


end behave;

