-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 15 19:22:35 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY AvanceFijo IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SI : IN STD_LOGIC := '0';
        SD : IN STD_LOGIC := '0';
        M0D : OUT STD_LOGIC;
        M1D : OUT STD_LOGIC;
        M0I : OUT STD_LOGIC;
        M1I : OUT STD_LOGIC
    );
END AvanceFijo;

ARCHITECTURE BEHAVIOR OF AvanceFijo IS
    TYPE type_fstate IS (Avanza_Recto,Corrige_Hacia_Derecha,Corrige_Hacia_Izquierda);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SI,SD)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Avanza_Recto;
            M0D <= '0';
            M1D <= '0';
            M0I <= '0';
            M1I <= '0';
        ELSE
            M0D <= '0';
            M1D <= '0';
            M0I <= '0';
            M1I <= '0';
            CASE fstate IS
                WHEN Avanza_Recto =>
                    IF (((SI = '1') AND (SD = '0'))) THEN
                        reg_fstate <= Corrige_Hacia_Derecha;
                    ELSIF (((SI = '0') AND (SD = '1'))) THEN
                        reg_fstate <= Corrige_Hacia_Izquierda;
                    ELSIF (((SI = '0') AND (SD = '0'))) THEN
                        reg_fstate <= Avanza_Recto;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Avanza_Recto;
                    END IF;

                    M0D <= '1';

                    M1D <= '0';

                    M0I <= '1';

                    M1I <= '0';
                WHEN Corrige_Hacia_Derecha =>
                    IF (((SI = '1') AND (SD = '0'))) THEN
                        reg_fstate <= Corrige_Hacia_Derecha;
                    ELSIF (((SI = '0') AND (SD = '0'))) THEN
                        reg_fstate <= Avanza_Recto;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Corrige_Hacia_Derecha;
                    END IF;

                    M0D <= '0';

                    M1D <= '1';

                    M0I <= '1';

                    M1I <= '0';
                WHEN Corrige_Hacia_Izquierda =>
                    IF (((SI = '0') AND (SD = '1'))) THEN
                        reg_fstate <= Corrige_Hacia_Izquierda;
                    ELSIF (((SI = '0') AND (SD = '0'))) THEN
                        reg_fstate <= Avanza_Recto;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Corrige_Hacia_Izquierda;
                    END IF;

                    M0D <= '1';

                    M1D <= '0';

                    M0I <= '0';

                    M1I <= '1';
                WHEN OTHERS => 
                    M0D <= 'X';
                    M1D <= 'X';
                    M0I <= 'X';
                    M1I <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
