LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TestADC is 

	port (
	CH1  : in std_logic_vector[11 downto 0];
	LED0 : out std_logic;
	LED1 : out std_logic
	);
	
end TestADC;

architecture behavioral of TestADC is

begin

	

end behavioral;
	