-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Nov 29 19:02:18 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY testBlock IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		w3 :  IN  STD_LOGIC;
		w10 :  IN  STD_LOGIC;
		w7 :  IN  STD_LOGIC;
		w0 :  IN  STD_LOGIC;
		w17 :  IN  STD_LOGIC;
		w21 :  IN  STD_LOGIC;
		w1 :  IN  STD_LOGIC;
		w4 :  IN  STD_LOGIC;
		w14 :  IN  STD_LOGIC;
		w11 :  IN  STD_LOGIC;
		w8 :  IN  STD_LOGIC;
		w22 :  IN  STD_LOGIC;
		w18 :  IN  STD_LOGIC;
		w15 :  IN  STD_LOGIC;
		w6 :  IN  STD_LOGIC;
		w2 :  IN  STD_LOGIC;
		w13 :  IN  STD_LOGIC;
		w9 :  IN  STD_LOGIC;
		w20 :  IN  STD_LOGIC;
		w16 :  IN  STD_LOGIC;
		w5 :  IN  STD_LOGIC;
		w12 :  IN  STD_LOGIC;
		w23 :  IN  STD_LOGIC;
		w19 :  IN  STD_LOGIC;
		Error :  OUT  STD_LOGIC;
		REG0_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG0_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG11_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG11_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG11_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG12_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG12_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG12_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG13_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG13_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG13_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG13_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG14_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG14_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG14_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG15_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG15_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG15_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG15_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG1_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG1_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG1_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG2_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG2_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG3_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG3_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG3_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG4_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG4_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG4_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG5_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG5_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG5_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG5_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG6_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG6_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG6_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG7_E :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG7_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG7_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG7_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG8_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG8_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG9_N :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG9_O :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG9_S :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END testBlock;

ARCHITECTURE bdf_type OF testBlock IS 

COMPONENT mux44
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT registrogenerico
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 RS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT d_ff
	PORT(D : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 Q : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT comparadorsumador4bit
	PORT(RegA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 RegB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 RegC : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 RegD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 RegOUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT vectorvalorcasilla
	PORT(		 int0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 int1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 int2 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 int3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 int4 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 int5 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 int6 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Vec_comp : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_231 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_232 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_233 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_234 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_235 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_236 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_237 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_238 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_240 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_241 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_242 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_243 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_244 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_245 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_246 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_247 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_248 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_249 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_250 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_251 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_252 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_253 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_254 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_255 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_256 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_257 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_258 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_259 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_260 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_261 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_262 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_263 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_264 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_265 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_266 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_267 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_268 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_269 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_270 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_271 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_272 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_273 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_274 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_275 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_276 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_277 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_278 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_279 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_280 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_281 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_282 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_283 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_284 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_164 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_170 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_172 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_285 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_286 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_287 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_182 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_183 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_184 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_288 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_191 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_192 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_289 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_198 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_199 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_290 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_206 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_208 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_209 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_210 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_211 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_218 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_219 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_291 :  STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN 
REG0_E <= SYNTHESIZED_WIRE_277;
REG0_S <= SYNTHESIZED_WIRE_276;
REG11_N <= SYNTHESIZED_WIRE_288;
REG11_O <= SYNTHESIZED_WIRE_192;
REG11_S <= SYNTHESIZED_WIRE_191;
REG12_E <= SYNTHESIZED_WIRE_198;
REG12_O <= SYNTHESIZED_WIRE_289;
REG12_S <= SYNTHESIZED_WIRE_199;
REG13_E <= SYNTHESIZED_WIRE_209;
REG13_N <= SYNTHESIZED_WIRE_210;
REG13_O <= SYNTHESIZED_WIRE_208;
REG13_S <= SYNTHESIZED_WIRE_211;
REG14_E <= SYNTHESIZED_WIRE_219;
REG14_N <= SYNTHESIZED_WIRE_291;
REG14_O <= SYNTHESIZED_WIRE_218;
REG15_E <= SYNTHESIZED_WIRE_10;
REG15_N <= SYNTHESIZED_WIRE_11;
REG15_O <= SYNTHESIZED_WIRE_9;
REG15_S <= SYNTHESIZED_WIRE_12;
REG1_E <= SYNTHESIZED_WIRE_83;
REG1_N <= SYNTHESIZED_WIRE_271;
REG1_S <= SYNTHESIZED_WIRE_82;
REG2_E <= SYNTHESIZED_WIRE_273;
REG2_N <= SYNTHESIZED_WIRE_272;
REG3_E <= SYNTHESIZED_WIRE_99;
REG3_N <= SYNTHESIZED_WIRE_274;
REG3_S <= SYNTHESIZED_WIRE_98;
REG4_E <= SYNTHESIZED_WIRE_278;
REG4_O <= SYNTHESIZED_WIRE_110;
REG4_S <= SYNTHESIZED_WIRE_111;
REG5_E <= SYNTHESIZED_WIRE_125;
REG5_N <= SYNTHESIZED_WIRE_123;
REG5_O <= SYNTHESIZED_WIRE_122;
REG5_S <= SYNTHESIZED_WIRE_124;
REG6_E <= SYNTHESIZED_WIRE_138;
REG6_N <= SYNTHESIZED_WIRE_137;
REG6_O <= SYNTHESIZED_WIRE_281;
REG7_E <= SYNTHESIZED_WIRE_172;
REG7_N <= SYNTHESIZED_WIRE_170;
REG7_O <= SYNTHESIZED_WIRE_169;
REG7_S <= SYNTHESIZED_WIRE_171;
REG8_O <= SYNTHESIZED_WIRE_286;
REG8_S <= SYNTHESIZED_WIRE_285;
REG9_N <= SYNTHESIZED_WIRE_287;
REG9_O <= SYNTHESIZED_WIRE_183;
REG9_S <= SYNTHESIZED_WIRE_182;



b2v_inst : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_231,
		 data0x => SYNTHESIZED_WIRE_232,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_276);


b2v_inst0 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_3,
		 RS => SYNTHESIZED_WIRE_4,
		 Q => SYNTHESIZED_WIRE_275);


b2v_inst1 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_5,
		 RS => SYNTHESIZED_WIRE_234,
		 Q => SYNTHESIZED_WIRE_232);


b2v_inst10 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_235,
		 RS => SYNTHESIZED_WIRE_235,
		 Q => SYNTHESIZED_WIRE_263);


b2v_inst100 : d_ff
PORT MAP(D => w19,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_240);


b2v_inst101 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_9,
		 RegB => SYNTHESIZED_WIRE_10,
		 RegC => SYNTHESIZED_WIRE_11,
		 RegD => SYNTHESIZED_WIRE_12,
		 RegOUT => SYNTHESIZED_WIRE_32);


b2v_inst102 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_236,
		 data0x => SYNTHESIZED_WIRE_237,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_10);


b2v_inst104 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_238,
		 data0x => SYNTHESIZED_WIRE_239,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_11);


b2v_inst105 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_240,
		 data0x => SYNTHESIZED_WIRE_241,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_12);


Error <= SYNTHESIZED_WIRE_242 AND SYNTHESIZED_WIRE_243;


b2v_inst11 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_24,
		 RS => SYNTHESIZED_WIRE_244,
		 Q => SYNTHESIZED_WIRE_237);


b2v_inst12 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_26,
		 RS => SYNTHESIZED_WIRE_245,
		 Q => SYNTHESIZED_WIRE_266);


b2v_inst13 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_28,
		 RS => SYNTHESIZED_WIRE_246,
		 Q => SYNTHESIZED_WIRE_239);


b2v_inst14 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_30,
		 RS => SYNTHESIZED_WIRE_244,
		 Q => SYNTHESIZED_WIRE_241);


b2v_inst15 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_32,
		 RS => SYNTHESIZED_WIRE_247,
		 Q => SYNTHESIZED_WIRE_270);


b2v_inst16 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_248,
		 data0x => SYNTHESIZED_WIRE_249,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_98);


b2v_inst17 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_250,
		 data0x => SYNTHESIZED_WIRE_251,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_82);


b2v_inst18 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_252,
		 data0x => SYNTHESIZED_WIRE_253,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_277);


b2v_inst19 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_254,
		 data0x => SYNTHESIZED_WIRE_255,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_83);


b2v_inst2 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_46,
		 RS => SYNTHESIZED_WIRE_246,
		 Q => SYNTHESIZED_WIRE_249);


b2v_inst20 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_256,
		 data0x => SYNTHESIZED_WIRE_257,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_273);


b2v_inst21 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_258,
		 data0x => SYNTHESIZED_WIRE_259,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_99);


b2v_inst22 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_260,
		 data0x => SYNTHESIZED_WIRE_261,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_287);


b2v_inst23 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_260,
		 data0x => SYNTHESIZED_WIRE_262,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_285);


b2v_inst24 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_242,
		 data0x => SYNTHESIZED_WIRE_263,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_191);


b2v_inst25 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_264,
		 data0x => SYNTHESIZED_WIRE_237,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_182);


b2v_inst26 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_265,
		 data0x => SYNTHESIZED_WIRE_266,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_278);


b2v_inst27 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_267,
		 data0x => SYNTHESIZED_WIRE_239,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_125);


b2v_inst28 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_268,
		 data0x => SYNTHESIZED_WIRE_241,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_138);


b2v_inst29 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_269,
		 data0x => SYNTHESIZED_WIRE_270,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_172);


b2v_inst3 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_78,
		 RS => SYNTHESIZED_WIRE_245,
		 Q => SYNTHESIZED_WIRE_251);


b2v_inst31 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_271,
		 RegB => SYNTHESIZED_WIRE_271,
		 RegC => SYNTHESIZED_WIRE_82,
		 RegD => SYNTHESIZED_WIRE_83,
		 RegOUT => SYNTHESIZED_WIRE_5);


b2v_inst32 : d_ff
PORT MAP(D => w3,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_231);


b2v_inst33 : d_ff
PORT MAP(D => w10,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_250);


b2v_inst34 : d_ff
PORT MAP(D => w7,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_254);


b2v_inst35 : d_ff
PORT MAP(D => w0,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_252);


b2v_inst36 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_272,
		 RegB => SYNTHESIZED_WIRE_272,
		 RegC => SYNTHESIZED_WIRE_273,
		 RegD => SYNTHESIZED_WIRE_273,
		 RegOUT => SYNTHESIZED_WIRE_46);


b2v_inst37 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_248,
		 data0x => SYNTHESIZED_WIRE_251,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_272);


b2v_inst38 : d_ff
PORT MAP(D => w17,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_248);


b2v_inst39 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_258,
		 data0x => SYNTHESIZED_WIRE_251,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_169);


b2v_inst4 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_94,
		 RS => SYNTHESIZED_WIRE_234,
		 Q => SYNTHESIZED_WIRE_253);


b2v_inst41 : d_ff
PORT MAP(D => w21,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_256);


b2v_inst42 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_274,
		 RegB => SYNTHESIZED_WIRE_274,
		 RegC => SYNTHESIZED_WIRE_98,
		 RegD => SYNTHESIZED_WIRE_99,
		 RegOUT => SYNTHESIZED_WIRE_78);


b2v_inst43 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_250,
		 data0x => SYNTHESIZED_WIRE_232,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_274);


b2v_inst45 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_252,
		 data0x => SYNTHESIZED_WIRE_275,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_110);


b2v_inst46 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_276,
		 RegB => SYNTHESIZED_WIRE_276,
		 RegC => SYNTHESIZED_WIRE_277,
		 RegD => SYNTHESIZED_WIRE_277,
		 RegOUT => SYNTHESIZED_WIRE_3);


b2v_inst47 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_110,
		 RegB => SYNTHESIZED_WIRE_111,
		 RegC => SYNTHESIZED_WIRE_278,
		 RegD => SYNTHESIZED_WIRE_278,
		 RegOUT => SYNTHESIZED_WIRE_94);


b2v_inst48 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_279,
		 data0x => SYNTHESIZED_WIRE_255,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_111);


b2v_inst49 : d_ff
PORT MAP(D => w4,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_279);


b2v_inst5 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_117,
		 RS => SYNTHESIZED_WIRE_245,
		 Q => SYNTHESIZED_WIRE_255);


b2v_inst50 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_254,
		 data0x => SYNTHESIZED_WIRE_232,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_122);


b2v_inst51 : d_ff
PORT MAP(D => w1,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_265);


b2v_inst52 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_122,
		 RegB => SYNTHESIZED_WIRE_123,
		 RegC => SYNTHESIZED_WIRE_124,
		 RegD => SYNTHESIZED_WIRE_125,
		 RegOUT => SYNTHESIZED_WIRE_117);


b2v_inst53 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_279,
		 data0x => SYNTHESIZED_WIRE_253,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_123);


b2v_inst54 : d_ff
PORT MAP(D => w14,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_258);


b2v_inst55 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_280,
		 data0x => SYNTHESIZED_WIRE_259,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_124);


b2v_inst555 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_231,
		 data0x => SYNTHESIZED_WIRE_275,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_271);


b2v_inst56 : d_ff
PORT MAP(D => w11,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_280);


b2v_inst57 : d_ff
PORT MAP(D => w8,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_267);


b2v_inst59 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_281,
		 RegB => SYNTHESIZED_WIRE_281,
		 RegC => SYNTHESIZED_WIRE_137,
		 RegD => SYNTHESIZED_WIRE_138,
		 RegOUT => SYNTHESIZED_WIRE_139);


b2v_inst6 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_139,
		 RS => SYNTHESIZED_WIRE_247,
		 Q => SYNTHESIZED_WIRE_257);


b2v_inst60 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_282,
		 data0x => SYNTHESIZED_WIRE_259,
		 result => SYNTHESIZED_WIRE_137);


b2v_inst61 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_256,
		 data0x => SYNTHESIZED_WIRE_249,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_281);


b2v_inst63 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_280,
		 data0x => SYNTHESIZED_WIRE_255,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_170);


b2v_inst64 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_267,
		 data0x => SYNTHESIZED_WIRE_255,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_208);


b2v_inst65 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_269,
		 data0x => SYNTHESIZED_WIRE_259,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_9);


b2v_inst67 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_283,
		 data0x => SYNTHESIZED_WIRE_261,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_198);


b2v_inst68 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_264,
		 data0x => SYNTHESIZED_WIRE_262,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_288);


b2v_inst69 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_284,
		 data0x => SYNTHESIZED_WIRE_262,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_209);


b2v_inst7 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_164,
		 RS => SYNTHESIZED_WIRE_246,
		 Q => SYNTHESIZED_WIRE_259);


b2v_inst70 : d_ff
PORT MAP(D => w18,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_282);


b2v_inst71 : d_ff
PORT MAP(D => w22,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_268);


b2v_inst72 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_282,
		 data0x => SYNTHESIZED_WIRE_257,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_171);


b2v_inst73 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_169,
		 RegB => SYNTHESIZED_WIRE_170,
		 RegC => SYNTHESIZED_WIRE_171,
		 RegD => SYNTHESIZED_WIRE_172,
		 RegOUT => SYNTHESIZED_WIRE_164);


b2v_inst74 : d_ff
PORT MAP(D => w15,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_269);


b2v_inst75 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_285,
		 RegB => SYNTHESIZED_WIRE_285,
		 RegC => SYNTHESIZED_WIRE_286,
		 RegD => SYNTHESIZED_WIRE_286,
		 RegOUT => SYNTHESIZED_WIRE_184);


b2v_inst76 : d_ff
PORT MAP(D => w6,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_260);


b2v_inst77 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_283,
		 data0x => SYNTHESIZED_WIRE_266,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_286);


b2v_inst78 : d_ff
PORT MAP(D => w2,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_283);


b2v_inst79 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_287,
		 RegB => SYNTHESIZED_WIRE_287,
		 RegC => SYNTHESIZED_WIRE_182,
		 RegD => SYNTHESIZED_WIRE_183,
		 RegOUT => SYNTHESIZED_WIRE_206);


b2v_inst8 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_184,
		 RS => SYNTHESIZED_WIRE_246,
		 Q => SYNTHESIZED_WIRE_261);


b2v_inst80 : d_ff
PORT MAP(D => w13,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_264);


b2v_inst81 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_284,
		 data0x => SYNTHESIZED_WIRE_239,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_183);


b2v_inst82 : d_ff
PORT MAP(D => w9,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_284);


b2v_inst83 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_288,
		 RegB => SYNTHESIZED_WIRE_288,
		 RegC => SYNTHESIZED_WIRE_191,
		 RegD => SYNTHESIZED_WIRE_192,
		 RegOUT => SYNTHESIZED_WIRE_24);


b2v_inst84 : d_ff
PORT MAP(D => w20,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_242);


b2v_inst85 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_236,
		 data0x => SYNTHESIZED_WIRE_270,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_192);


b2v_inst86 : d_ff
PORT MAP(D => w16,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_236);


b2v_inst87 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_289,
		 RegB => SYNTHESIZED_WIRE_289,
		 RegC => SYNTHESIZED_WIRE_198,
		 RegD => SYNTHESIZED_WIRE_199,
		 RegOUT => SYNTHESIZED_WIRE_26);


b2v_inst88 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_265,
		 data0x => SYNTHESIZED_WIRE_253,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_289);


b2v_inst89 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_290,
		 data0x => SYNTHESIZED_WIRE_239,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_199);


b2v_inst9 : registrogenerico
PORT MAP(clk => clk,
		 reset => reset,
		 D => SYNTHESIZED_WIRE_206,
		 RS => SYNTHESIZED_WIRE_247,
		 Q => SYNTHESIZED_WIRE_262);


b2v_inst90 : d_ff
PORT MAP(D => w5,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_290);


b2v_inst91 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_208,
		 RegB => SYNTHESIZED_WIRE_209,
		 RegC => SYNTHESIZED_WIRE_210,
		 RegD => SYNTHESIZED_WIRE_211,
		 RegOUT => SYNTHESIZED_WIRE_28);


b2v_inst92 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_290,
		 data0x => SYNTHESIZED_WIRE_266,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_210);


b2v_inst93 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_238,
		 data0x => SYNTHESIZED_WIRE_270,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_211);


b2v_inst94 : d_ff
PORT MAP(D => w12,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_238);


b2v_inst95 : comparadorsumador4bit
PORT MAP(RegA => SYNTHESIZED_WIRE_218,
		 RegB => SYNTHESIZED_WIRE_219,
		 RegC => SYNTHESIZED_WIRE_291,
		 RegD => SYNTHESIZED_WIRE_291,
		 RegOUT => SYNTHESIZED_WIRE_30);


b2v_inst96 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_268,
		 data0x => SYNTHESIZED_WIRE_257,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_218);


b2v_inst97 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_243,
		 data0x => SYNTHESIZED_WIRE_263,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_219);


b2v_inst98 : d_ff
PORT MAP(D => w23,
		 clk => clk,
		 reset => reset,
		 Q => SYNTHESIZED_WIRE_243);


b2v_inst99 : mux44
PORT MAP(sel => SYNTHESIZED_WIRE_240,
		 data0x => SYNTHESIZED_WIRE_270,
		 data1x => SYNTHESIZED_WIRE_233,
		 result => SYNTHESIZED_WIRE_291);


b2v_instvecval : vectorvalorcasilla
PORT MAP(		 int0 => SYNTHESIZED_WIRE_235,
		 int1 => SYNTHESIZED_WIRE_244,
		 int2 => SYNTHESIZED_WIRE_247,
		 int3 => SYNTHESIZED_WIRE_246,
		 int4 => SYNTHESIZED_WIRE_245,
		 int5 => SYNTHESIZED_WIRE_234,
		 int6 => SYNTHESIZED_WIRE_4,
		 Vec_comp => SYNTHESIZED_WIRE_233);


END bdf_type;